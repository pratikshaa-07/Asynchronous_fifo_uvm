package fifo_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "define.sv"
  `include "wrt_seq_item.sv"
  `include "rd_seq_item.sv"

  `include "wrt_sequence.sv"
  `include "rd_sequence.sv"

  `include "write_sequencer.sv"
  `include "read_sequencer.sv"

  `include "write_driver.sv"
  `include "read_driver.sv"

  `include "write_mon.sv"
  `include "read_mon.sv"

  `include "write_agent.sv"
  `include "read_agent.sv"

  `include "subscriber.sv"
  `include "scoreboard.sv"

  `include "virtual_sequencer.sv"
  `include "virtual_sequence.sv"

  `include "environment.sv"
  `include "test.sv"

endpackage

